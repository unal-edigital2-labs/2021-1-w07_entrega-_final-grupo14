`timescale 1ns / 1ps

module infrarrojo(
  input [4:0] infras,
  output [4:0] infras2
);

  assign infras2 = infras;

endmodule